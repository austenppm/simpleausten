module externalIn(input [15:0] in,
				output [15:0] mdr_inputSource);
	assign mdr_inputSource = in ;	
endmodule
						